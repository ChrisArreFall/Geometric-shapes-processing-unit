module draw #(parameter N)
				(input logic [N-1:0] x, y, xc, yc
				 output logic [N*8:0] s);
	//x = a
	//y = b
	//xc = c
	//yc = d
	logic C0,C1,C2,C3,C4,C5,C6,C7;
	assign C0 = 
	initial begin
	//si es circulo o elipse entonces 
    s = {};
	end
	assign s[] = a | b; // OR
	
	x*N+y
endmodule